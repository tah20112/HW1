// Simple program to print hello
module hello_test();
initial begin
	$display("Hello, CompArch!");
end
endmodule
